module clock_counter(
	input logic clk_in,
	output logic clk_out
);

//insert clock module here

endmodule