module mux2( 	input logic [15:0] keyboard_data, button_ 
				input logic [15:0] button_data,
				input logic sel,
				output logic [15:0] SNES_data);
