module clk_counter(
input logic clk_i,
output logic clk_slow
);

//write clock divider here

endmodule