/***************************************
* Affiliation: Oregon State University
* Author: Cody McCall
*
* Course: ECE 271 - Digital Logic Design
* Project Name: ECE 271 Design Project
* Team Number: 09
*
* Description: Ps2 Keyboard Top Module
* Start Date: 06/03/2018
*
****************************************/
module ps2_Top(
input logic ps2_data, clk_15khz,
output logic [15:0] ps2_data);

	
endmodule 